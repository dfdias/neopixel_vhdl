NeoPixel_receiver.vhd

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity NeoPixel_receiver is --this module will receive some data from serial port
port()
end NeoPixel_receiver;

architecture Behav of NeoPixel_receiver is
signal
